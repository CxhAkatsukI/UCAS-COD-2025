// timescale directive: simulation time unit is 10ns, precision is 1ns
`timescale 10ns / 1ns

// Macro definitions for bus widths
`define ADDR_WIDTH 5  // Register file address width
`define DATA_WIDTH 32 // Data bus width

//==============================================================================
// Module: simple_cpu
// Description: A simple MIPS-like CPU core with integrated control logic.
//              (Code organized by strict pipeline stage definitions)
//==============================================================================
module simple_cpu (
    //-- Global Signals --
    input         clk,            // Clock signal
    input         rst,            // Reset signal

    //-- Instruction Fetch Interface --
    output [31:0] PC,             // Program Counter output
    input  [31:0] Instruction,    // Instruction input from memory

    //-- Data Memory Interface --
    output [31:0] Address,        // Memory address output
    output        MemWrite,       // Memory write enable signal
    output [31:0] Write_data,     // Data to write to memory
    output [ 3:0] Write_strb,     // Memory byte strobes for writes
    input  [31:0] Read_data,      // Data read from memory
    output        MemRead         // Memory read enable signal
);

  //----------------------------------------------------------------------------
  // Internal Wires - Connecting Logic Blocks and Modules
  // (Grouped here for clarity, used across stages)
  //----------------------------------------------------------------------------

  //-- Signals generated in ID (purely from Instruction) --
  wire [ 5:0] opcode;               // Opcode field
  wire [ 4:0] rs;                   // Source register 1 specifier
  wire [ 4:0] rt;                   // Source register 2 specifier / Branch Func
  wire [ 4:0] rd;                   // Destination register specifier (R-type)
  wire [ 4:0] shamt;                // Shift amount (R-type shift)
  wire [ 5:0] funct;                // Function field (R-type)
  wire [15:0] imm_16;               // 16-bit immediate value
  wire [25:0] imm_J;                // 26-bit immediate for jump
  wire [31:0] imm_SE;               // Sign-extended immediate
  wire [31:0] imm_0E;               // Zero-extended immediate
  wire [31:0] imm_B_ext;            // Sign-extended branch immediate
  wire [31:0] lui_result;           // Result for LUI instruction
  wire        use_zero_extend;      // Control for immediate extension type
  reg  [ 4:0] current_state;        // Current state of the FSM
  reg  [ 4:0] next_state;           // Next state of the FSM
  reg  [31:0] IR;                   // Instruction Register (holds current instruction)

  wire        reg_dst_input;          // Selects destination register (rd/rt/ra hint)
  wire        is_branch;              // Indicates Branch instruction
  wire        branch_condition_satisfied; // Indicates branch condition is satisfied
  wire        mem_read_internal;      // Internal Memory read enable (Load)
  wire        mem_write_internal;     // Internal Memory write enable (Store)
  wire        alu_src_imm_input;      // Selects ALU source 2 (Reg/Imm)
  wire        reg_write_cond;         // Precondition for register write enable (base check)
  wire        alu_op_ok;              // Indicates ALUOp can be derived from opcode
  wire [ 2:0] alu_op_cond;            // ALU operation hint from opcode
  wire        is_alu_operation;       // Indicates an ALU operation is needed
  wire        is_shift_operation;     // Indicates a Shift operation is needed
  wire [ 2:0] alu_op;                 // Decoded ALU operation (R/I type)
  wire [ 1:0] shifter_op;             // Decoded Shift operation type
  wire        is_shamt;               // Indicates shamt is used for shift amount
  wire        is_zero_cmp;            // Indicates branch compares rs against zero
  wire        is_move;                // Indicates MOVZ/MOVN
  wire        is_lui;                 // Indicates LUI instruction
  wire        is_load_store;          // Indicates Load/Store instruction
  wire [ 2:0] move_alu_op;            // ALU operation code for MOVZ/MOVN
  wire        is_jump;                // Indicates any Jump instruction occurred (J, JAL, JR, JALR)
  wire        is_link_jump;           // Indicates JAL or JALR instruction
  wire        is_j_instr;
  wire        is_jal_instr;
  wire        is_jr_instr;
  wire        is_jalr_instr;
  wire        is_REGIMM;
  wire        NOP;                    // Indicates NOP instruction (all bits 0)
  wire        write_disallowed;       // Instr. type that never writes back
  wire        intermediate_reg_write_cond; // Base write condition refined

  //-- Signals from Register File (ID Stage Read) --
  wire [31:0] RF_rdata1;              // Data read from RegFile port 1 (rs)
  wire [31:0] RF_rdata2;              // Data read from RegFile port 2 (rt)

  //-- Signals from/for PC Path (Generated/Used across stages) --
  wire [31:0] next_pc;                // Next program counter value (Calculated in EX)
  wire [31:0] current_pc;             // Current program counter value (from PC module in IF)
  wire [31:0] pc_store;               // PC+8 for JAL/JALR link address (Calculated in EX)

  //-- Signals from ALU/Shifter Path (Generated in EX) --
  wire [31:0] alu_src1;               // First ALU operand
  wire [31:0] alu_src2;               // Second ALU operand
  wire [31:0] shifter_src1;           // First Shifter operand (data)
  wire [31:0] shifter_src2;           // Second Shifter operand (shift amount)
  wire [ 2:0] alu_op_final;           // Final ALU operation control to ALU
  wire        alu_zero;               // ALU Zero flag
  reg  [31:0] alu_result;             // ALU computation result
  reg  [31:0] shift_result;           // Shifter result

  //-- Signals from Memory Path (Generated in MEM) --
  wire [31:0] load_data;              // Data processed from memory/registers for load operations

  //-- Signals for WB Stage --
  wire        RF_wen;                 // Final write enable to RegFile
  wire [ 4:0] RF_waddr;               // Write address to RegFile
  reg  [31:0] RF_wdata;               // Write data to RegFile


  //============================================================================
  // PIPELINE STAGE 0: FSM Implementation
  //============================================================================

  // -- FSM State Definitions --
  localparam IF = 5'b00001,
             ID = 5'b00010,
             EX = 5'b00100,
             MEM = 5'b01000,
             WB = 5'b10000;

  // -- FSM State Register --
  always @(posedge clk) begin
    if (rst) begin
      current_state <= IF;         // Reset state
    end else begin
      current_state <= next_state; // Update state based on FSM logic
    end
  end

  // -- FSM Next State Logic --
  always @(*) begin
    case (current_state)
      IF : next_state = ID;
      ID : begin
            if (NOP) begin
              next_state = IF;
            end
            else begin
              next_state = EX;
            end
      end
      EX : begin
        if (is_j_instr || is_REGIMM || is_branch) begin
          next_state = IF;
        end
        else if (is_load_store) begin
          next_state = MEM;
        end
        else begin
          next_state = WB;
        end
      end
      MEM : begin
        if (opcode[3]) begin
          next_state = IF;
        end
        else begin
          next_state = WB;
        end
      end
      WB : next_state = IF;
      default: next_state = IF;
  endcase
  end

  // -- FSM Output Logic --
  assign IRWrite = current_state[0];
  assign Regwrite_fsm = current_state[4];

  // -- Instruction Register Logic --
  always @(posedge clk) begin
    if (IRWrite) begin
      IR <= Instruction; // Reset instruction register
    end else begin
      IR <= IR;          // Fetch instruction from memory
    end
  end


  //============================================================================
  // PIPELINE STAGE 1: Instruction Fetch (IF)
  //============================================================================

  //-- PC Register --
  wire pc_write_enable = (current_state == IF) ||                                          // Always update after IF (for PC+4 usually)
                       ((current_state == EX) && is_jump) ||                               // Update for any jump in EX
                       ((current_state == EX) && is_branch && branch_condition_satisfied); // Update for taken branch in EX
  pc instance_pc (
      .clk        (clk),
      .rst        (rst),
      .pc_write_enable (pc_write_enable), // Input: PC write enable signal (from control logic)
      .next_pc    (next_pc),              // Input: Next PC value (Calculated in EX stage)
      .pc         (current_pc)            // Output: Current PC value (Used across stages)
  );


  //============================================================================
  // PIPELINE STAGE 2: Instruction Decode / Register Fetch (ID)
  //============================================================================

  //-- Instruction Field Decoding --
  assign      opcode   = IR[31:26]; // Opcode field
  assign      rs       = IR[25:21]; // Source register 1 specifier
  assign      rt       = IR[20:16]; // Source register 2 specifier / Branch Func
  assign      rd       = IR[15:11]; // Destination register specifier (R-type)
  assign      shamt    = IR[10: 6]; // Shift amount (R-type shift)
  assign      funct    = IR[ 5: 0]; // Function field (R-type)
  assign      imm_16   = IR[15: 0]; // 16-bit immediate value
  assign      imm_J    = IR[25: 0]; // 26-bit immediate for jump

  //-- Immediate Value Processing (Purely from Instruction) --
  assign      NOP      = (~|IR);                                      // NOP instruction (all bits 0)
  assign      imm_SE   = {{16{imm_16[15]}}, imm_16};                  // Sign-extended immediate
  assign      imm_0E   = {16'b0, imm_16};                             // Zero-extended immediate
  assign      imm_B_ext= {{16{imm_16[15]}}, imm_16};                  // Sign-extended branch immediate (used in EX)
  assign      lui_result = {imm_16, 16'b0};                           // Result for LUI instruction (used in WB)
  assign      use_zero_extend = (opcode[5:3] == 3'b001) && opcode[2]; // Use Zero Ext for ANDI/ORI/XORI (used in EX)

  //-- Primary Control Signal Generation (Purely from Instruction) --
  wire        is_branch_sub     = (opcode[5:2] == 4'b0001);                    // Specific branch types
  wire        is_branch_slt     = (opcode == 6'b000001);                       // Branches that use slt as alu_op
  assign      is_branch         = (is_branch_sub || is_branch_slt);            // General branch flag
  assign      reg_dst_input     = opcode[5] ^ opcode[3];                       // Hint for WB Stage dest reg sel
  assign      mem_read_internal = current_state[3] && (opcode[5:3] == 3'b100); // Control for MEM Stage
  assign      mem_write_internal= current_state[3] && (opcode[5:3] == 3'b101); // Control for MEM Stage
  assign      alu_src_imm_input = ((opcode[5] || opcode[3]) && !opcode[4]);    // Control for EX Stage (ALU Src Sel)

  //-- Secondary Control Signal Generation (Purely from Instruction or derived ID signals) --
  wire        imm_arithmetic    = (opcode[5:3] == 3'b001 && ~&opcode[2:0]);       // I-type Arith?
  assign      is_load_store     = opcode[5:3] == 3'b100 || opcode[5:3] == 3'b101; // Load or Store?
  assign      reg_write_cond    = !mem_write_internal && !is_branch;              // Base RegWrite condition (used in WB)

  // -- Decode I-type arith op based on opcode --
  wire [ 2:0] arith_type;
  assign      arith_type[0]     = (~opcode[2] & opcode[1]) | (opcode[2] & opcode[0]);
  assign      arith_type[1]     = ~opcode[2];
  assign      arith_type[2]     = opcode[1] & ~opcode[0];
  assign      alu_op_cond       = is_branch_slt  ? 3'b111 :
                                  is_branch_sub  ? 3'b110 :
                                  is_load_store  ? 3'b010 :
                                  imm_arithmetic ? arith_type :
                                  3'bxxx;
  assign      alu_op_ok         = (imm_arithmetic || is_branch || is_load_store);      // Validity of hint for EX

  assign      is_alu_operation   = ((~|opcode && funct[5] == 1'b1) || imm_arithmetic); // Is it an ALU op? (Used EX/WB)
  assign      is_shift_operation = (~|opcode && ~|funct[5:3]);                         // Is it a Shift op? (Used EX/WB)

  // -- Decode R-type arith op based on funct --
  wire [ 2:0] r_type_arith_op;
  assign      r_type_arith_op[0] = (funct[3] & funct[1]) | (~funct[3] & funct[2] & funct[0]);
  assign      r_type_arith_op[1] = funct[3] | ~funct[2];
  assign      r_type_arith_op[2] = (funct[3] & ~funct[0]) | (~funct[3] & funct[1]);
  assign      alu_op             = (~|opcode) ? r_type_arith_op : alu_op_cond ;        // Base ALU op (R/I type) (Used EX)

  // -- Decode R-type shift op based on funct --
  wire [ 1:0] shift_type;                                                              // Decode R-type shift op based on funct
  assign      shift_type[0]      = funct[1] & funct[0];
  assign      shift_type[1]      = funct[1];
  assign      shifter_op         = is_shift_operation ? shift_type : 2'b00;            // Shift op type (Used EX)
  assign      is_shamt           = is_shift_operation && ~funct[2];                    // Use shamt? (Used EX)

  assign      is_zero_cmp        = is_branch && (opcode[2:0] == 3'b110 || opcode[2:0] == 3'b111 || opcode[2:0] == 3'b001); // Compare rs to 0? (Used EX)

  assign      is_move            = (~|opcode && funct[1] && funct[3] && !funct[5]);    // MOVZ/MOVN? (Used EX/WB)
  assign      is_lui             = (opcode == 6'b001111);                              // LUI? (Used WB)
  assign      move_alu_op        = 3'b001;                                             // ALU Op for Move (Used EX)

  assign      is_j_instr         = (opcode == 6'b000010);
  assign      is_jal_instr       = (opcode == 6'b000011);
  assign      is_jr_instr        = (~|opcode && funct == 6'b001000);
  assign      is_jalr_instr      = (~|opcode && funct == 6'b001001);
  assign      is_jump            = is_j_instr || is_jal_instr || is_jr_instr || is_jalr_instr; // Is it any Jump? (Used EX)
  assign      is_link_jump       = is_jal_instr || is_jalr_instr;                              // Is it JAL/JALR? (Used EX/WB)
  assign      is_REGIMM          = (opcode == 6'b000001);                                      // Is it REGIMM? (Used EX)

  assign      write_disallowed   = is_j_instr || is_jr_instr || mem_write_internal;            // Instr. that don't write back (refined) (Used WB)
  assign      intermediate_reg_write_cond = reg_write_cond && !write_disallowed;               // Base write condition refined (Used WB)




  //-- Register File Read --
  reg_file instance_reg_file (
      .clk        (clk),
      .waddr      (RF_waddr),         // Input: Write address (From WB stage)
      .raddr1     (rs),               // Input: Read address 1 (rs field from ID)
      .raddr2     (rt),               // Input: Read address 2 (rt field from ID)
      .wen        (RF_wen),           // Input: Write enable (From WB stage)
      .wdata      (RF_wdata),         // Input: Write data (From WB stage)
      .rdata1     (RF_rdata1),        // Output: Read data 1 (rs value) -> To EX
      .rdata2     (RF_rdata2)         // Output: Read data 2 (rt value) -> To EX/MEM/WB
  );

  //============================================================================
  // PIPELINE STAGE 3: Execute (EX)
  //============================================================================

  //-- ALU Source Selector Logic (Uses ID signals, Reg Data) --
  assign      alu_src1           = (is_move) ? 32'b0 : RF_rdata1;                         // ALU Input A
  assign      alu_src2           = (is_zero_cmp)       ? 32'b0 :                          // ALU Input B
                                   (alu_src_imm_input) ? (use_zero_extend ? imm_0E : imm_SE) :
                                   RF_rdata2;

  //-- Shifter Source Selector Logic (Uses ID signals, Reg Data) --
  assign      shifter_src1       = RF_rdata2;                                             // Shifter Input A (Data)
  assign      shifter_src2       = (is_shamt) ? {27'b0, shamt} : {27'b0, RF_rdata1[4:0]}; // Shifter Input B (Amount)

  //-- ALU Op Generator Logic (Uses ID signals) --
  assign      alu_op_final       = (is_move)          ? move_alu_op :
                                   (is_alu_operation) ? alu_op :
                                   (alu_op_ok)        ? alu_op_cond :
                                   3'b010;                                                // Final ALU Op -> To ALU

  //-- ALU Execution --
  wire [31:0] alu_out;                // ALU computation result

  alu instance_alu (
      .A          (alu_src1),         // Input A from Src Sel
      .B          (alu_src2),         // Input B from Src Sel
      .ALUop      (alu_op_final),     // Input Opcode from Op Gen
      .Overflow   (),
      .CarryOut   (),
      .Zero       (alu_zero),         // Output: Zero flag -> To EX (PC Ctrl), WB
      .Result     (alu_out)           // Output: ALU computation result -> To EX (PC Ctrl), MEM, WB
  );

  always @(posedge clk) begin
      alu_result <= alu_out;          // Store ALU result for MEM stage
  end

  //-- Shifter Execution --
  wire [31:0] shifter_out;                // Shifter computation result

  shifter instance_shifter (
      .A          (shifter_src1),         // Input Data from Src Sel
      .B          (shifter_src2[4:0]),    // Input Shift Amount from Src Sel
      .Shiftop    (shifter_op),           // Input Opcode from ID
      .Result     (shifter_out)           // Output: Shifter result -> To WB
  );

  always @(posedge clk) begin
      shift_result <= shifter_out;        // Store Shifter result for WB stage
  end

  //-- PC Controller Logic (Uses ID signals, EX results, IF PC) --
  assign      branch_condition_satisfied = is_branch &&                                                                    // Check using signals from ID and results from EX
                                           ( (is_branch_slt && (rt[0] ^ alu_result[0])) ||                                 // REGIMM check using rt(funct_branch) from ID, alu_result from EX
                                             (is_branch_sub && opcode[1] && (opcode[0] ^ (alu_result[31] || alu_zero))) || // BLEZ/BGTZ check using opcode from ID, alu_result/zero from EX
                                             (is_branch_sub && !opcode[1] && (opcode[0] ^ alu_zero))                       // BEQ/BNE check using opcode from ID, alu_zero from EX
                                           );

  wire [31:0] branch_target      = (current_pc) + (imm_B_ext << 2);                                                   // Branch target addr calculation

  wire [31:0] jump_target        = (is_j_instr || is_jal_instr) ? {current_pc[31:28], imm_J, 2'b00} : RF_rdata1;      // J/JAL or JR/JALR target calculation

  // Next PC Selection based on control signals (ID) and conditions (EX)
  assign      next_pc            = (rst)                                                    ? 32'h00000000 :          // Reset PC value
                                   (current_state == EX && is_jump)                         ? jump_target  :          // Jump target selection
                                   (current_state == EX && is_branch && branch_condition_satisfied) ? branch_target : // Branch target selection
                                   current_pc + 4;                                                                    // Default: PC + 4 -> To IF

  // PC+8 Calculation for Link Instructions (Uses ID signal, IF PC)
  assign      pc_store           = is_link_jump ? (current_pc + 4) : 32'b0;                                           // Value to store for JAL/JALR -> To WB

  //============================================================================
  // PIPELINE STAGE 4: Memory Access (MEM)
  //============================================================================

  //-- Load/Store Address and Data Logic (Uses ID signals, EX results, ID reg data) --
  wire [ 1:0] addr_offset        = alu_result[1:0];            // Byte offset (from EX result)
  wire        addr_0             = (addr_offset == 2'b00);
  wire        addr_1             = (addr_offset == 2'b01);
  wire        addr_2             = (addr_offset == 2'b10);
  wire        addr_3             = (addr_offset == 2'b11);

  // Memory Address Output Calculation (Uses EX result)
  assign      Address            = {alu_result[31:2], 2'b00};  // Word-aligned address -> To Memory Interface

  // Memory Write Strobe Generation (Uses ID signals, EX result offset)
  assign      Write_strb         = {4{mem_write_internal}} & ( // Use is_store (mem_write_internal) from ID
                                     (({4{opcode[1:0] == 2'b00}} & ((addr_0 ? 4'b0001 : 0) | (addr_1 ? 4'b0010 : 0) | (addr_2 ? 4'b0100 : 0) | (addr_3 ? 4'b1000 : 0))) | // SB
                                     ({4{opcode[1:0] == 2'b01}} & ((addr_0 ? 4'b0011 : 0) | (addr_2 ? 4'b1100 : 0))) |                                                    // SH
                                     ({4{opcode[1:0] == 2'b11}} & (addr_0 ? 4'b1111 : 4'b0000)) |                                                                         // SW
                                     ({4{opcode[2:0] == 3'b010}} & ((addr_0 ? 4'b0001 : 0) | (addr_1 ? 4'b0011 : 0) | (addr_2 ? 4'b0111 : 0) | (addr_3 ? 4'b1111 : 0))) | // SWL
                                     ({4{opcode[2:0] == 3'b110}} & ((addr_0 ? 4'b1111 : 0) | (addr_1 ? 4'b1110 : 0) | (addr_2 ? 4'b1100 : 0) | (addr_3 ? 4'b1000 : 0)))   // SWR
                                    )); // -> To Memory Interface

  assign      Write_data         = {32{mem_write_internal}} & ( // Format RF_rdata2 for stores -> To Memory Interface
                                     (({32{opcode[1:0] == 2'b00}} & {4{RF_rdata2[7:0]}}) | // SB
                                     ({32{opcode[1:0] == 2'b01}} & {2{RF_rdata2[15:0]}}) | // SH
                                     ({32{opcode[1:0] == 2'b11}} & RF_rdata2) |            // SW
                                     ({32{opcode[2:0] == 3'b010}} & ( // SWL (Logic kept as-is)
                                         (addr_0 ? {24'b0, RF_rdata2[31:24]} :
                                          addr_1 ? {16'b0, RF_rdata2[31:16]} :
                                          addr_2 ? { 8'b0, RF_rdata2[31: 8]} :
                                                   RF_rdata2)
                                     )) |
                                     ({32{opcode[2:0] == 3'b110}} & ( // SWR (Logic kept as-is)
                                         (addr_0 ? RF_rdata2 :
                                          addr_1 ? {RF_rdata2[23:0],  8'b0} :
                                          addr_2 ? {RF_rdata2[15:0], 16'b0} :
                                                   {RF_rdata2[ 7:0], 24'b0})
                                     )))
                                   );

   // Processing of Data Read from Memory (Uses ID signals, EX result offset, ID reg data, Mem input)
   assign      load_data          = mem_read_internal ? // Process Read_data -> To WB Stage
                                    ( (opcode[1:0] == 2'b00) ?  // LB/LBU
                                      (addr_0 ? {{24{(~opcode[2] & Read_data [ 7])}}, Read_data [ 7: 0]} :
                                       addr_1 ? {{24{(~opcode[2] & Read_data [15])}}, Read_data [15: 8]} :
                                       addr_2 ? {{24{(~opcode[2] & Read_data [23])}}, Read_data [23:16]} :
                                                {{24{(~opcode[2] & Read_data [31])}}, Read_data [31:24]} )

                                    : (opcode[1:0] == 2'b01) ?  // LH/LHU
                                      (addr_0 ? {{16{(~opcode[2] & Read_data [15])}}, Read_data [15: 0]} :
                                       addr_2 ? {{16{(~opcode[2] & Read_data [31])}}, Read_data [31:16]} :
                                                32'b0 )

                                    : (opcode[1:0] == 2'b11) ? Read_data // LW

                                    : (opcode[2:0] == 3'b010) ? // LWL
                                      (addr_0 ? {Read_data [ 7: 0], RF_rdata2 [23: 0]} :
                                       addr_1 ? {Read_data [15: 0], RF_rdata2 [15: 0]} :
                                       addr_2 ? {Read_data [23: 0], RF_rdata2 [ 7: 0]} :
                                                Read_data )

                                    : (opcode[2:0] == 3'b110) ? // LWR
                                      (addr_0 ? Read_data :
                                       addr_1 ? {RF_rdata2 [31:24], Read_data [31: 8]} :
                                       addr_2 ? {RF_rdata2 [31:16], Read_data [31:16]} :
                                                {RF_rdata2 [31: 8], Read_data [31:24]} )

                                    : 32'b0 ) // Default unknown load
                                    : 32'b0;  // Default if not a load


  //============================================================================
  // PIPELINE STAGE 5: Write Back (WB)
  //============================================================================

  //-- Register Write Address and Enable Logic (Uses ID signals, EX results) --
  assign      RF_waddr           = (is_link_jump) ? 5'd31 :           // JAL/JALR -> $ra (from ID)
                                   (reg_dst_input) ? rt :             // I-type/Load hint -> rt (from ID)
                                   rd;                                // R-type hint -> rd (from ID)
                                                                      // -> To RegFile instance

  assign      RF_wen             = Regwrite_fsm & ((intermediate_reg_write_cond && !is_move) || // Use conditions from ID and...
                                   (is_move && (funct[0] ^ alu_zero) && reg_write_cond));       // ...MOVZ/N check using alu_zero from EX
                                                                                                // -> To RegFile instance

  //-- Write Back Data Selection (Uses ID signals, EX results, MEM results) --
  wire [31:0] _RF_wdata;                                                       // Write data to RegFile (processed from ID, EX, MEM)
  assign      _RF_wdata          = (is_lui)             ? lui_result :         // P1: LUI (from ID)
                                   (mem_read_internal)  ? load_data :          // P2: Load result from MEM
                                   (is_move)            ? RF_rdata1 :          // P3: MOVZ/MOVN result (rs) from ID
                                   (is_alu_operation)   ? alu_result :         // P4: Other ALU result from EX
                                   (is_shift_operation) ? shift_result :       // P5: Shifter result from EX
                                   (is_link_jump)       ? pc_store :           // P6: Link address (PC+8) from EX
                                   32'b0;                                      // Default: 0 (No writeback)
                                                                               // -> To RegFile instance
  always @(posedge clk) begin
      RF_wdata <= _RF_wdata;                                                   // Store write data for RegFile
  end

  //----------------------------------------------------------------------------
  // Top-Level Output Assignments
  //----------------------------------------------------------------------------
  assign      PC                 = current_pc;                      // Output current PC (from IF stage)
  assign      MemWrite           = mem_write_internal;              // Output MemWrite signal (from ID stage control)
  assign      MemRead            = mem_read_internal;               // Output MemRead signal (from ID stage control)

endmodule


//==============================================================================
// Module: pc (Remains unchanged)
// Description: Program Counter register. Stores the address of the next
//              instruction to be fetched.
//==============================================================================
module pc (
    input         clk,
    input         rst,
    input         pc_write_enable,
    input  [31:0] next_pc,
    output reg [31:0] pc
);
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      pc <= 32'h00000000;
    end else if (pc_write_enable) begin
      pc <= next_pc;
    end
  end
endmodule

